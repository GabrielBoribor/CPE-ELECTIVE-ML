module Full_Decoder(a1,a2,a3,b1,b2,b3,b4,b5,b6,b7);
input a1,a2,a3;
output b1,b2,b3,b4,b5,b6,b7;
endmodule