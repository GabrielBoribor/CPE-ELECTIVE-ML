module test_and(a1,a2,b);
input a1,a2;
output b;

endmodule