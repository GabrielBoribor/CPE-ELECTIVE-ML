module Decoder(a1,a2,b1,b2,b3);
input a1,a2;
output b1,b2,b3;
endmodule