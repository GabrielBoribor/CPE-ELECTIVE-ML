module test_nor(a1,a2,b);
input a1,a2;
output b;

endmodule