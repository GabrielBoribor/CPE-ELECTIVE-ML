module test_not(a1,b);
input a1;
output b;

endmodule